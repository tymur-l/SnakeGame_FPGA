`ifndef init_vh
`define init_vh

`include "./define.vh"

`define GRID_INIT game_grid[0][0] = 4'b1100;\
game_grid[0][1] = 4'b1100;\
game_grid[0][2] = 4'b1100;\
game_grid[0][3] = 4'b1100;\
game_grid[0][4] = 4'b1100;\
game_grid[0][5] = 4'b1100;\
game_grid[0][6] = 4'b1100;\
game_grid[0][7] = 4'b1100;\
game_grid[0][8] = 4'b1100;\
game_grid[0][9] = 4'b1100;\
game_grid[0][10] = 4'b1100;\
game_grid[0][11] = 4'b1100;\
game_grid[0][12] = 4'b1100;\
game_grid[0][13] = 4'b1100;\
game_grid[0][14] = 4'b1100;\
game_grid[0][15] = 4'b1100;\
game_grid[0][16] = 4'b1100;\
game_grid[0][17] = 4'b1100;\
game_grid[0][18] = 4'b1100;\
game_grid[0][19] = 4'b1100;\
game_grid[0][20] = 4'b1100;\
game_grid[0][21] = 4'b1100;\
game_grid[0][22] = 4'b1100;\
game_grid[0][23] = 4'b1100;\
game_grid[0][24] = 4'b1100;\
game_grid[0][25] = 4'b1100;\
game_grid[0][26] = 4'b1100;\
game_grid[0][27] = 4'b1100;\
game_grid[0][28] = 4'b1100;\
game_grid[0][29] = 4'b1100;\
game_grid[1][0] = 4'b1100;\
game_grid[1][1] = 4'b1100;\
game_grid[1][2] = 4'b1100;\
game_grid[1][3] = 4'b1100;\
game_grid[1][4] = 4'b1100;\
game_grid[1][5] = 4'b1100;\
game_grid[1][6] = 4'b1100;\
game_grid[1][7] = 4'b1100;\
game_grid[1][8] = 4'b1100;\
game_grid[1][9] = 4'b1100;\
game_grid[1][10] = 4'b1100;\
game_grid[1][11] = 4'b1100;\
game_grid[1][12] = 4'b1100;\
game_grid[1][13] = 4'b1100;\
game_grid[1][14] = 4'b1100;\
game_grid[1][15] = 4'b1100;\
game_grid[1][16] = 4'b1100;\
game_grid[1][17] = 4'b1100;\
game_grid[1][18] = 4'b1100;\
game_grid[1][19] = 4'b1100;\
game_grid[1][20] = 4'b1100;\
game_grid[1][21] = 4'b1100;\
game_grid[1][22] = 4'b1100;\
game_grid[1][23] = 4'b1100;\
game_grid[1][24] = 4'b1100;\
game_grid[1][25] = 4'b1100;\
game_grid[1][26] = 4'b1100;\
game_grid[1][27] = 4'b1100;\
game_grid[1][28] = 4'b1100;\
game_grid[1][29] = 4'b1100;\
game_grid[2][0] = 4'b1100;\
game_grid[2][1] = 4'b1100;\
game_grid[2][2] = 4'b1100;\
game_grid[2][3] = 4'b1100;\
game_grid[2][4] = 4'b1100;\
game_grid[2][5] = 4'b1100;\
game_grid[2][6] = 4'b1100;\
game_grid[2][7] = 4'b1100;\
game_grid[2][8] = 4'b1100;\
game_grid[2][9] = 4'b1100;\
game_grid[2][10] = 4'b1100;\
game_grid[2][11] = 4'b1100;\
game_grid[2][12] = 4'b1100;\
game_grid[2][13] = 4'b1100;\
game_grid[2][14] = 4'b1100;\
game_grid[2][15] = 4'b1100;\
game_grid[2][16] = 4'b1100;\
game_grid[2][17] = 4'b1100;\
game_grid[2][18] = 4'b1100;\
game_grid[2][19] = 4'b1100;\
game_grid[2][20] = 4'b1100;\
game_grid[2][21] = 4'b1100;\
game_grid[2][22] = 4'b1100;\
game_grid[2][23] = 4'b1100;\
game_grid[2][24] = 4'b1100;\
game_grid[2][25] = 4'b1100;\
game_grid[2][26] = 4'b1100;\
game_grid[2][27] = 4'b1100;\
game_grid[2][28] = 4'b1100;\
game_grid[2][29] = 4'b1100;\
game_grid[3][0] = 4'b1100;\
game_grid[3][1] = 4'b1100;\
game_grid[3][2] = 4'b1100;\
game_grid[3][3] = 4'b1100;\
game_grid[3][4] = 4'b1100;\
game_grid[3][5] = 4'b1100;\
game_grid[3][6] = 4'b1100;\
game_grid[3][7] = 4'b1100;\
game_grid[3][8] = 4'b1100;\
game_grid[3][9] = 4'b1100;\
game_grid[3][10] = 4'b1100;\
game_grid[3][11] = 4'b1100;\
game_grid[3][12] = 4'b1100;\
game_grid[3][13] = 4'b1100;\
game_grid[3][14] = 4'b1100;\
game_grid[3][15] = 4'b1100;\
game_grid[3][16] = 4'b1100;\
game_grid[3][17] = 4'b1100;\
game_grid[3][18] = 4'b1100;\
game_grid[3][19] = 4'b1100;\
game_grid[3][20] = 4'b1100;\
game_grid[3][21] = 4'b1100;\
game_grid[3][22] = 4'b1100;\
game_grid[3][23] = 4'b1100;\
game_grid[3][24] = 4'b1100;\
game_grid[3][25] = 4'b1100;\
game_grid[3][26] = 4'b1100;\
game_grid[3][27] = 4'b1100;\
game_grid[3][28] = 4'b1100;\
game_grid[3][29] = 4'b1100;\
game_grid[4][0] = 4'b1100;\
game_grid[4][1] = 4'b1100;\
game_grid[4][2] = 4'b1100;\
game_grid[4][3] = 4'b1100;\
game_grid[4][4] = 4'b1100;\
game_grid[4][5] = 4'b1100;\
game_grid[4][6] = 4'b1100;\
game_grid[4][7] = 4'b1100;\
game_grid[4][8] = 4'b1100;\
game_grid[4][9] = 4'b1100;\
game_grid[4][10] = 4'b1100;\
game_grid[4][11] = 4'b1100;\
game_grid[4][12] = 4'b1100;\
game_grid[4][13] = 4'b1100;\
game_grid[4][14] = 4'b1100;\
game_grid[4][15] = 4'b1100;\
game_grid[4][16] = 4'b1100;\
game_grid[4][17] = 4'b1100;\
game_grid[4][18] = 4'b1100;\
game_grid[4][19] = 4'b1100;\
game_grid[4][20] = 4'b1100;\
game_grid[4][21] = 4'b1100;\
game_grid[4][22] = 4'b1100;\
game_grid[4][23] = 4'b1100;\
game_grid[4][24] = 4'b1100;\
game_grid[4][25] = 4'b1100;\
game_grid[4][26] = 4'b1100;\
game_grid[4][27] = 4'b1100;\
game_grid[4][28] = 4'b1100;\
game_grid[4][29] = 4'b1100;\
game_grid[5][0] = 4'b1100;\
game_grid[5][1] = 4'b1100;\
game_grid[5][2] = 4'b1100;\
game_grid[5][3] = 4'b1100;\
game_grid[5][4] = 4'b1100;\
game_grid[5][5] = 4'b1100;\
game_grid[5][6] = 4'b1100;\
game_grid[5][7] = 4'b1100;\
game_grid[5][8] = 4'b1100;\
game_grid[5][9] = 4'b1100;\
game_grid[5][10] = 4'b1100;\
game_grid[5][11] = 4'b1100;\
game_grid[5][12] = 4'b1100;\
game_grid[5][13] = 4'b1100;\
game_grid[5][14] = 4'b1100;\
game_grid[5][15] = 4'b1100;\
game_grid[5][16] = 4'b1100;\
game_grid[5][17] = 4'b1100;\
game_grid[5][18] = 4'b1100;\
game_grid[5][19] = 4'b1100;\
game_grid[5][20] = 4'b1100;\
game_grid[5][21] = 4'b1100;\
game_grid[5][22] = 4'b1100;\
game_grid[5][23] = 4'b1100;\
game_grid[5][24] = 4'b1100;\
game_grid[5][25] = 4'b1100;\
game_grid[5][26] = 4'b1100;\
game_grid[5][27] = 4'b1100;\
game_grid[5][28] = 4'b1100;\
game_grid[5][29] = 4'b1100;\
game_grid[6][0] = 4'b1100;\
game_grid[6][1] = 4'b1100;\
game_grid[6][2] = 4'b1100;\
game_grid[6][3] = 4'b1100;\
game_grid[6][4] = 4'b1100;\
game_grid[6][5] = 4'b1100;\
game_grid[6][6] = 4'b1100;\
game_grid[6][7] = 4'b1100;\
game_grid[6][8] = 4'b1100;\
game_grid[6][9] = 4'b1100;\
game_grid[6][10] = 4'b1100;\
game_grid[6][11] = 4'b1100;\
game_grid[6][12] = 4'b1100;\
game_grid[6][13] = 4'b1100;\
game_grid[6][14] = 4'b1100;\
game_grid[6][15] = 4'b1100;\
game_grid[6][16] = 4'b1100;\
game_grid[6][17] = 4'b1100;\
game_grid[6][18] = 4'b1100;\
game_grid[6][19] = 4'b1100;\
game_grid[6][20] = 4'b1100;\
game_grid[6][21] = 4'b1100;\
game_grid[6][22] = 4'b1100;\
game_grid[6][23] = 4'b1100;\
game_grid[6][24] = 4'b1100;\
game_grid[6][25] = 4'b1100;\
game_grid[6][26] = 4'b1100;\
game_grid[6][27] = 4'b1100;\
game_grid[6][28] = 4'b1100;\
game_grid[6][29] = 4'b1100;\
game_grid[7][0] = 4'b1100;\
game_grid[7][1] = 4'b1100;\
game_grid[7][2] = 4'b1100;\
game_grid[7][3] = 4'b1100;\
game_grid[7][4] = 4'b1100;\
game_grid[7][5] = 4'b1100;\
game_grid[7][6] = 4'b1100;\
game_grid[7][7] = 4'b1100;\
game_grid[7][8] = 4'b1100;\
game_grid[7][9] = 4'b1100;\
game_grid[7][10] = 4'b1100;\
game_grid[7][11] = 4'b1100;\
game_grid[7][12] = 4'b1100;\
game_grid[7][13] = 4'b1100;\
game_grid[7][14] = 4'b1100;\
game_grid[7][15] = 4'b1100;\
game_grid[7][16] = 4'b1100;\
game_grid[7][17] = 4'b1100;\
game_grid[7][18] = 4'b1100;\
game_grid[7][19] = 4'b1100;\
game_grid[7][20] = 4'b1100;\
game_grid[7][21] = 4'b1100;\
game_grid[7][22] = 4'b1100;\
game_grid[7][23] = 4'b1100;\
game_grid[7][24] = 4'b1100;\
game_grid[7][25] = 4'b1100;\
game_grid[7][26] = 4'b1100;\
game_grid[7][27] = 4'b1100;\
game_grid[7][28] = 4'b1100;\
game_grid[7][29] = 4'b1100;\
game_grid[8][0] = 4'b1100;\
game_grid[8][1] = 4'b1100;\
game_grid[8][2] = 4'b1100;\
game_grid[8][3] = 4'b1100;\
game_grid[8][4] = 4'b1100;\
game_grid[8][5] = 4'b1100;\
game_grid[8][6] = 4'b1100;\
game_grid[8][7] = 4'b1100;\
game_grid[8][8] = 4'b1100;\
game_grid[8][9] = 4'b1100;\
game_grid[8][10] = 4'b1100;\
game_grid[8][11] = 4'b1100;\
game_grid[8][12] = 4'b1100;\
game_grid[8][13] = 4'b1100;\
game_grid[8][14] = 4'b1100;\
game_grid[8][15] = 4'b1100;\
game_grid[8][16] = 4'b1100;\
game_grid[8][17] = 4'b1100;\
game_grid[8][18] = 4'b1100;\
game_grid[8][19] = 4'b1100;\
game_grid[8][20] = 4'b1100;\
game_grid[8][21] = 4'b1100;\
game_grid[8][22] = 4'b1100;\
game_grid[8][23] = 4'b1100;\
game_grid[8][24] = 4'b1100;\
game_grid[8][25] = 4'b1100;\
game_grid[8][26] = 4'b1100;\
game_grid[8][27] = 4'b1100;\
game_grid[8][28] = 4'b1100;\
game_grid[8][29] = 4'b1100;\
game_grid[9][0] = 4'b1100;\
game_grid[9][1] = 4'b1100;\
game_grid[9][2] = 4'b1100;\
game_grid[9][3] = 4'b1100;\
game_grid[9][4] = 4'b1100;\
game_grid[9][5] = 4'b1100;\
game_grid[9][6] = 4'b1100;\
game_grid[9][7] = 4'b1100;\
game_grid[9][8] = 4'b1100;\
game_grid[9][9] = 4'b1100;\
game_grid[9][10] = 4'b1100;\
game_grid[9][11] = 4'b1100;\
game_grid[9][12] = 4'b1100;\
game_grid[9][13] = 4'b1100;\
game_grid[9][14] = 4'b1100;\
game_grid[9][15] = 4'b1100;\
game_grid[9][16] = 4'b1100;\
game_grid[9][17] = 4'b1100;\
game_grid[9][18] = 4'b1100;\
game_grid[9][19] = 4'b1100;\
game_grid[9][20] = 4'b1100;\
game_grid[9][21] = 4'b1100;\
game_grid[9][22] = 4'b1100;\
game_grid[9][23] = 4'b1100;\
game_grid[9][24] = 4'b1100;\
game_grid[9][25] = 4'b1100;\
game_grid[9][26] = 4'b1100;\
game_grid[9][27] = 4'b1100;\
game_grid[9][28] = 4'b1100;\
game_grid[9][29] = 4'b1100;\
game_grid[10][0] = 4'b1100;\
game_grid[10][1] = 4'b1100;\
game_grid[10][2] = 4'b1100;\
game_grid[10][3] = 4'b1100;\
game_grid[10][4] = 4'b1100;\
game_grid[10][5] = 4'b1100;\
game_grid[10][6] = 4'b1100;\
game_grid[10][7] = 4'b1100;\
game_grid[10][8] = 4'b1100;\
game_grid[10][9] = 4'b1100;\
game_grid[10][10] = 4'b1100;\
game_grid[10][11] = 4'b1100;\
game_grid[10][12] = 4'b1100;\
game_grid[10][13] = 4'b1100;\
game_grid[10][14] = 4'b1100;\
game_grid[10][15] = 4'b1100;\
game_grid[10][16] = 4'b1100;\
game_grid[10][17] = 4'b1100;\
game_grid[10][18] = 4'b1100;\
game_grid[10][19] = 4'b1100;\
game_grid[10][20] = 4'b1100;\
game_grid[10][21] = 4'b1100;\
game_grid[10][22] = 4'b1100;\
game_grid[10][23] = 4'b1100;\
game_grid[10][24] = 4'b1100;\
game_grid[10][25] = 4'b1100;\
game_grid[10][26] = 4'b1100;\
game_grid[10][27] = 4'b1100;\
game_grid[10][28] = 4'b1100;\
game_grid[10][29] = 4'b1100;\
game_grid[11][0] = 4'b1100;\
game_grid[11][1] = 4'b1100;\
game_grid[11][2] = 4'b1100;\
game_grid[11][3] = 4'b1100;\
game_grid[11][4] = 4'b1100;\
game_grid[11][5] = 4'b1100;\
game_grid[11][6] = 4'b1100;\
game_grid[11][7] = 4'b1100;\
game_grid[11][8] = 4'b1100;\
game_grid[11][9] = 4'b1100;\
game_grid[11][10] = 4'b1100;\
game_grid[11][11] = 4'b1100;\
game_grid[11][12] = 4'b1100;\
game_grid[11][13] = 4'b1100;\
game_grid[11][14] = 4'b1100;\
game_grid[11][15] = 4'b1100;\
game_grid[11][16] = 4'b1100;\
game_grid[11][17] = 4'b1100;\
game_grid[11][18] = 4'b1100;\
game_grid[11][19] = 4'b1100;\
game_grid[11][20] = 4'b1100;\
game_grid[11][21] = 4'b1100;\
game_grid[11][22] = 4'b1100;\
game_grid[11][23] = 4'b1100;\
game_grid[11][24] = 4'b1100;\
game_grid[11][25] = 4'b1100;\
game_grid[11][26] = 4'b1100;\
game_grid[11][27] = 4'b1100;\
game_grid[11][28] = 4'b1100;\
game_grid[11][29] = 4'b1100;\
game_grid[12][0] = 4'b1100;\
game_grid[12][1] = 4'b1100;\
game_grid[12][2] = 4'b1100;\
game_grid[12][3] = 4'b1100;\
game_grid[12][4] = 4'b1100;\
game_grid[12][5] = 4'b1100;\
game_grid[12][6] = 4'b1100;\
game_grid[12][7] = 4'b1100;\
game_grid[12][8] = 4'b1100;\
game_grid[12][9] = 4'b1100;\
game_grid[12][10] = 4'b1100;\
game_grid[12][11] = 4'b1100;\
game_grid[12][12] = 4'b1100;\
game_grid[12][13] = 4'b1100;\
game_grid[12][14] = 4'b1100;\
game_grid[12][15] = 4'b1100;\
game_grid[12][16] = 4'b1100;\
game_grid[12][17] = 4'b1100;\
game_grid[12][18] = 4'b1100;\
game_grid[12][19] = 4'b1100;\
game_grid[12][20] = 4'b1100;\
game_grid[12][21] = 4'b1100;\
game_grid[12][22] = 4'b1100;\
game_grid[12][23] = 4'b1100;\
game_grid[12][24] = 4'b1100;\
game_grid[12][25] = 4'b1100;\
game_grid[12][26] = 4'b1100;\
game_grid[12][27] = 4'b1100;\
game_grid[12][28] = 4'b1100;\
game_grid[12][29] = 4'b1100;\
game_grid[13][0] = 4'b1100;\
game_grid[13][1] = 4'b1100;\
game_grid[13][2] = 4'b1100;\
game_grid[13][3] = 4'b1100;\
game_grid[13][4] = 4'b1100;\
game_grid[13][5] = 4'b1100;\
game_grid[13][6] = 4'b1100;\
game_grid[13][7] = 4'b1100;\
game_grid[13][8] = 4'b1100;\
game_grid[13][9] = 4'b1100;\
game_grid[13][10] = 4'b1100;\
game_grid[13][11] = 4'b1100;\
game_grid[13][12] = 4'b1100;\
game_grid[13][13] = 4'b1100;\
game_grid[13][14] = 4'b1100;\
game_grid[13][15] = 4'b1100;\
game_grid[13][16] = 4'b1100;\
game_grid[13][17] = 4'b1100;\
game_grid[13][18] = 4'b1100;\
game_grid[13][19] = 4'b1100;\
game_grid[13][20] = 4'b1100;\
game_grid[13][21] = 4'b1100;\
game_grid[13][22] = 4'b1100;\
game_grid[13][23] = 4'b1100;\
game_grid[13][24] = 4'b1100;\
game_grid[13][25] = 4'b1100;\
game_grid[13][26] = 4'b1100;\
game_grid[13][27] = 4'b1100;\
game_grid[13][28] = 4'b1100;\
game_grid[13][29] = 4'b1100;\
game_grid[14][0] = 4'b1100;\
game_grid[14][1] = 4'b1100;\
game_grid[14][2] = 4'b1100;\
game_grid[14][3] = 4'b1100;\
game_grid[14][4] = 4'b1100;\
game_grid[14][5] = 4'b1100;\
game_grid[14][6] = 4'b1100;\
game_grid[14][7] = 4'b1100;\
game_grid[14][8] = 4'b1100;\
game_grid[14][9] = 4'b1100;\
game_grid[14][10] = 4'b1100;\
game_grid[14][11] = 4'b1100;\
game_grid[14][12] = 4'b1100;\
game_grid[14][13] = 4'b1100;\
game_grid[14][14] = 4'b1100;\
game_grid[14][15] = 4'b1100;\
game_grid[14][16] = 4'b1100;\
game_grid[14][17] = 4'b1100;\
game_grid[14][18] = 4'b1100;\
game_grid[14][19] = 4'b1100;\
game_grid[14][20] = 4'b1100;\
game_grid[14][21] = 4'b1100;\
game_grid[14][22] = 4'b1100;\
game_grid[14][23] = 4'b1100;\
game_grid[14][24] = 4'b1100;\
game_grid[14][25] = 4'b1100;\
game_grid[14][26] = 4'b1100;\
game_grid[14][27] = 4'b1100;\
game_grid[14][28] = 4'b1100;\
game_grid[14][29] = 4'b1100;\
game_grid[15][0] = 4'b1100;\
game_grid[15][1] = 4'b1100;\
game_grid[15][2] = 4'b1100;\
game_grid[15][3] = 4'b1100;\
game_grid[15][4] = 4'b1100;\
game_grid[15][5] = 4'b1100;\
game_grid[15][6] = 4'b1100;\
game_grid[15][7] = 4'b1100;\
game_grid[15][8] = 4'b1100;\
game_grid[15][9] = 4'b1100;\
game_grid[15][10] = 4'b1100;\
game_grid[15][11] = 4'b1100;\
game_grid[15][12] = 4'b1100;\
game_grid[15][13] = 4'b1100;\
game_grid[15][14] = 4'b1100;\
game_grid[15][15] = 4'b1100;\
game_grid[15][16] = 4'b1100;\
game_grid[15][17] = 4'b1100;\
game_grid[15][18] = 4'b1100;\
game_grid[15][19] = 4'b1100;\
game_grid[15][20] = 4'b1100;\
game_grid[15][21] = 4'b1100;\
game_grid[15][22] = 4'b1100;\
game_grid[15][23] = 4'b1100;\
game_grid[15][24] = 4'b1100;\
game_grid[15][25] = 4'b1100;\
game_grid[15][26] = 4'b1100;\
game_grid[15][27] = 4'b1100;\
game_grid[15][28] = 4'b1100;\
game_grid[15][29] = 4'b1100;\
game_grid[16][0] = 4'b1100;\
game_grid[16][1] = 4'b1100;\
game_grid[16][2] = 4'b1100;\
game_grid[16][3] = 4'b1100;\
game_grid[16][4] = 4'b1100;\
game_grid[16][5] = 4'b1100;\
game_grid[16][6] = 4'b1100;\
game_grid[16][7] = 4'b1100;\
game_grid[16][8] = 4'b1100;\
game_grid[16][9] = 4'b1100;\
game_grid[16][10] = 4'b1100;\
game_grid[16][11] = 4'b1100;\
game_grid[16][12] = 4'b1100;\
game_grid[16][13] = 4'b1100;\
game_grid[16][14] = 4'b1100;\
game_grid[16][15] = 4'b1100;\
game_grid[16][16] = 4'b1100;\
game_grid[16][17] = 4'b1100;\
game_grid[16][18] = 4'b1100;\
game_grid[16][19] = 4'b1100;\
game_grid[16][20] = 4'b1100;\
game_grid[16][21] = 4'b1100;\
game_grid[16][22] = 4'b1100;\
game_grid[16][23] = 4'b1100;\
game_grid[16][24] = 4'b1100;\
game_grid[16][25] = 4'b1100;\
game_grid[16][26] = 4'b1100;\
game_grid[16][27] = 4'b1100;\
game_grid[16][28] = 4'b1100;\
game_grid[16][29] = 4'b1100;\
game_grid[17][0] = 4'b1100;\
game_grid[17][1] = 4'b1100;\
game_grid[17][2] = 4'b1100;\
game_grid[17][3] = 4'b1100;\
game_grid[17][4] = 4'b1100;\
game_grid[17][5] = 4'b1100;\
game_grid[17][6] = 4'b1100;\
game_grid[17][7] = 4'b1100;\
game_grid[17][8] = 4'b1100;\
game_grid[17][9] = 4'b1100;\
game_grid[17][10] = 4'b1100;\
game_grid[17][11] = 4'b1100;\
game_grid[17][12] = 4'b1100;\
game_grid[17][13] = 4'b1100;\
game_grid[17][14] = 4'b1100;\
game_grid[17][15] = 4'b1100;\
game_grid[17][16] = 4'b1100;\
game_grid[17][17] = 4'b1100;\
game_grid[17][18] = 4'b1100;\
game_grid[17][19] = 4'b1100;\
game_grid[17][20] = 4'b1100;\
game_grid[17][21] = 4'b1100;\
game_grid[17][22] = 4'b1100;\
game_grid[17][23] = 4'b1100;\
game_grid[17][24] = 4'b1100;\
game_grid[17][25] = 4'b1100;\
game_grid[17][26] = 4'b1100;\
game_grid[17][27] = 4'b1100;\
game_grid[17][28] = 4'b1100;\
game_grid[17][29] = 4'b1100;\
game_grid[18][0] = 4'b1100;\
game_grid[18][1] = 4'b1100;\
game_grid[18][2] = 4'b1100;\
game_grid[18][3] = 4'b1100;\
game_grid[18][4] = 4'b1100;\
game_grid[18][5] = 4'b1100;\
game_grid[18][6] = 4'b1100;\
game_grid[18][7] = 4'b1100;\
game_grid[18][8] = 4'b1100;\
game_grid[18][9] = 4'b1100;\
game_grid[18][10] = 4'b1100;\
game_grid[18][11] = 4'b1100;\
game_grid[18][12] = 4'b1100;\
game_grid[18][13] = 4'b1100;\
game_grid[18][14] = 4'b1100;\
game_grid[18][15] = 4'b1100;\
game_grid[18][16] = 4'b1100;\
game_grid[18][17] = 4'b1100;\
game_grid[18][18] = 4'b1100;\
game_grid[18][19] = 4'b1100;\
game_grid[18][20] = 4'b1100;\
game_grid[18][21] = 4'b1100;\
game_grid[18][22] = 4'b1100;\
game_grid[18][23] = 4'b1100;\
game_grid[18][24] = 4'b1100;\
game_grid[18][25] = 4'b1100;\
game_grid[18][26] = 4'b1100;\
game_grid[18][27] = 4'b1100;\
game_grid[18][28] = 4'b1100;\
game_grid[18][29] = 4'b1100;\
game_grid[19][0] = 4'b1100;\
game_grid[19][1] = 4'b1100;\
game_grid[19][2] = 4'b1100;\
game_grid[19][3] = 4'b1100;\
game_grid[19][4] = 4'b1100;\
game_grid[19][5] = 4'b1100;\
game_grid[19][6] = 4'b1100;\
game_grid[19][7] = 4'b1100;\
game_grid[19][8] = 4'b1100;\
game_grid[19][9] = 4'b1100;\
game_grid[19][10] = 4'b1100;\
game_grid[19][11] = 4'b1100;\
game_grid[19][12] = 4'b1100;\
game_grid[19][13] = 4'b1100;\
game_grid[19][14] = {`ENT_SNAKE_HEAD, 2'b00};\
game_grid[19][15] = 4'b1100;\
game_grid[19][16] = 4'b1100;\
game_grid[19][17] = 4'b1100;\
game_grid[19][18] = 4'b1100;\
game_grid[19][19] = 4'b1100;\
game_grid[19][20] = 4'b1100;\
game_grid[19][21] = 4'b1100;\
game_grid[19][22] = 4'b1100;\
game_grid[19][23] = 4'b1100;\
game_grid[19][24] = 4'b1100;\
game_grid[19][25] = 4'b1100;\
game_grid[19][26] = 4'b1100;\
game_grid[19][27] = 4'b1100;\
game_grid[19][28] = 4'b1100;\
game_grid[19][29] = 4'b1100;\
game_grid[20][0] = 4'b1100;\
game_grid[20][1] = 4'b1100;\
game_grid[20][2] = 4'b1100;\
game_grid[20][3] = 4'b1100;\
game_grid[20][4] = 4'b1100;\
game_grid[20][5] = 4'b1100;\
game_grid[20][6] = 4'b1100;\
game_grid[20][7] = 4'b1100;\
game_grid[20][8] = 4'b1100;\
game_grid[20][9] = 4'b1100;\
game_grid[20][10] = 4'b1100;\
game_grid[20][11] = 4'b1100;\
game_grid[20][12] = 4'b1100;\
game_grid[20][13] = 4'b1100;\
game_grid[20][14] = 4'b1100;\
game_grid[20][15] = 4'b1100;\
game_grid[20][16] = 4'b1100;\
game_grid[20][17] = 4'b1100;\
game_grid[20][18] = 4'b1100;\
game_grid[20][19] = 4'b1100;\
game_grid[20][20] = 4'b1100;\
game_grid[20][21] = 4'b1100;\
game_grid[20][22] = 4'b1100;\
game_grid[20][23] = 4'b1100;\
game_grid[20][24] = 4'b1100;\
game_grid[20][25] = 4'b1100;\
game_grid[20][26] = 4'b1100;\
game_grid[20][27] = 4'b1100;\
game_grid[20][28] = 4'b1100;\
game_grid[20][29] = 4'b1100;\
game_grid[21][0] = 4'b1100;\
game_grid[21][1] = 4'b1100;\
game_grid[21][2] = 4'b1100;\
game_grid[21][3] = 4'b1100;\
game_grid[21][4] = 4'b1100;\
game_grid[21][5] = 4'b1100;\
game_grid[21][6] = 4'b1100;\
game_grid[21][7] = 4'b1100;\
game_grid[21][8] = 4'b1100;\
game_grid[21][9] = 4'b1100;\
game_grid[21][10] = 4'b1100;\
game_grid[21][11] = 4'b1100;\
game_grid[21][12] = 4'b1100;\
game_grid[21][13] = 4'b1100;\
game_grid[21][14] = 4'b1100;\
game_grid[21][15] = 4'b1100;\
game_grid[21][16] = 4'b1100;\
game_grid[21][17] = 4'b1100;\
game_grid[21][18] = 4'b1100;\
game_grid[21][19] = 4'b1100;\
game_grid[21][20] = 4'b1100;\
game_grid[21][21] = 4'b1100;\
game_grid[21][22] = 4'b1100;\
game_grid[21][23] = 4'b1100;\
game_grid[21][24] = 4'b1100;\
game_grid[21][25] = 4'b1100;\
game_grid[21][26] = 4'b1100;\
game_grid[21][27] = 4'b1100;\
game_grid[21][28] = 4'b1100;\
game_grid[21][29] = 4'b1100;\
game_grid[22][0] = 4'b1100;\
game_grid[22][1] = 4'b1100;\
game_grid[22][2] = 4'b1100;\
game_grid[22][3] = 4'b1100;\
game_grid[22][4] = 4'b1100;\
game_grid[22][5] = 4'b1100;\
game_grid[22][6] = 4'b1100;\
game_grid[22][7] = 4'b1100;\
game_grid[22][8] = 4'b1100;\
game_grid[22][9] = 4'b1100;\
game_grid[22][10] = 4'b1100;\
game_grid[22][11] = 4'b1100;\
game_grid[22][12] = 4'b1100;\
game_grid[22][13] = 4'b1100;\
game_grid[22][14] = 4'b1100;\
game_grid[22][15] = 4'b1100;\
game_grid[22][16] = 4'b1100;\
game_grid[22][17] = 4'b1100;\
game_grid[22][18] = 4'b1100;\
game_grid[22][19] = 4'b1100;\
game_grid[22][20] = 4'b1100;\
game_grid[22][21] = 4'b1100;\
game_grid[22][22] = 4'b1100;\
game_grid[22][23] = 4'b1100;\
game_grid[22][24] = 4'b1100;\
game_grid[22][25] = 4'b1100;\
game_grid[22][26] = 4'b1100;\
game_grid[22][27] = 4'b1100;\
game_grid[22][28] = 4'b1100;\
game_grid[22][29] = 4'b1100;\
game_grid[23][0] = 4'b1100;\
game_grid[23][1] = 4'b1100;\
game_grid[23][2] = 4'b1100;\
game_grid[23][3] = 4'b1100;\
game_grid[23][4] = 4'b1100;\
game_grid[23][5] = 4'b1100;\
game_grid[23][6] = 4'b1100;\
game_grid[23][7] = 4'b1100;\
game_grid[23][8] = 4'b1100;\
game_grid[23][9] = 4'b1100;\
game_grid[23][10] = 4'b1100;\
game_grid[23][11] = 4'b1100;\
game_grid[23][12] = 4'b1100;\
game_grid[23][13] = 4'b1100;\
game_grid[23][14] = 4'b1100;\
game_grid[23][15] = 4'b1100;\
game_grid[23][16] = 4'b1100;\
game_grid[23][17] = 4'b1100;\
game_grid[23][18] = 4'b1100;\
game_grid[23][19] = 4'b1100;\
game_grid[23][20] = 4'b1100;\
game_grid[23][21] = 4'b1100;\
game_grid[23][22] = 4'b1100;\
game_grid[23][23] = 4'b1100;\
game_grid[23][24] = 4'b1100;\
game_grid[23][25] = 4'b1100;\
game_grid[23][26] = 4'b1100;\
game_grid[23][27] = 4'b1100;\
game_grid[23][28] = 4'b1100;\
game_grid[23][29] = 4'b1100;\
game_grid[24][0] = 4'b1100;\
game_grid[24][1] = 4'b1100;\
game_grid[24][2] = 4'b1100;\
game_grid[24][3] = 4'b1100;\
game_grid[24][4] = 4'b1100;\
game_grid[24][5] = 4'b1100;\
game_grid[24][6] = 4'b1100;\
game_grid[24][7] = 4'b1100;\
game_grid[24][8] = 4'b1100;\
game_grid[24][9] = 4'b1100;\
game_grid[24][10] = 4'b1100;\
game_grid[24][11] = 4'b1100;\
game_grid[24][12] = 4'b1100;\
game_grid[24][13] = 4'b1100;\
game_grid[24][14] = 4'b1100;\
game_grid[24][15] = 4'b1100;\
game_grid[24][16] = 4'b1100;\
game_grid[24][17] = 4'b1100;\
game_grid[24][18] = 4'b1100;\
game_grid[24][19] = 4'b1100;\
game_grid[24][20] = 4'b1100;\
game_grid[24][21] = 4'b1100;\
game_grid[24][22] = 4'b1100;\
game_grid[24][23] = 4'b1100;\
game_grid[24][24] = 4'b1100;\
game_grid[24][25] = 4'b1100;\
game_grid[24][26] = 4'b1100;\
game_grid[24][27] = 4'b1100;\
game_grid[24][28] = 4'b1100;\
game_grid[24][29] = 4'b1100;\
game_grid[25][0] = 4'b1100;\
game_grid[25][1] = 4'b1100;\
game_grid[25][2] = 4'b1100;\
game_grid[25][3] = 4'b1100;\
game_grid[25][4] = 4'b1100;\
game_grid[25][5] = 4'b1100;\
game_grid[25][6] = 4'b1100;\
game_grid[25][7] = 4'b1100;\
game_grid[25][8] = 4'b1100;\
game_grid[25][9] = 4'b1100;\
game_grid[25][10] = 4'b1100;\
game_grid[25][11] = 4'b1100;\
game_grid[25][12] = 4'b1100;\
game_grid[25][13] = 4'b1100;\
game_grid[25][14] = 4'b1100;\
game_grid[25][15] = 4'b1100;\
game_grid[25][16] = 4'b1100;\
game_grid[25][17] = 4'b1100;\
game_grid[25][18] = 4'b1100;\
game_grid[25][19] = 4'b1100;\
game_grid[25][20] = 4'b1100;\
game_grid[25][21] = 4'b1100;\
game_grid[25][22] = 4'b1100;\
game_grid[25][23] = 4'b1100;\
game_grid[25][24] = 4'b1100;\
game_grid[25][25] = 4'b1100;\
game_grid[25][26] = 4'b1100;\
game_grid[25][27] = 4'b1100;\
game_grid[25][28] = 4'b1100;\
game_grid[25][29] = 4'b1100;\
game_grid[26][0] = 4'b1100;\
game_grid[26][1] = 4'b1100;\
game_grid[26][2] = 4'b1100;\
game_grid[26][3] = 4'b1100;\
game_grid[26][4] = 4'b1100;\
game_grid[26][5] = 4'b1100;\
game_grid[26][6] = 4'b1100;\
game_grid[26][7] = 4'b1100;\
game_grid[26][8] = 4'b1100;\
game_grid[26][9] = 4'b1100;\
game_grid[26][10] = 4'b1100;\
game_grid[26][11] = 4'b1100;\
game_grid[26][12] = 4'b1100;\
game_grid[26][13] = 4'b1100;\
game_grid[26][14] = 4'b1100;\
game_grid[26][15] = 4'b1100;\
game_grid[26][16] = 4'b1100;\
game_grid[26][17] = 4'b1100;\
game_grid[26][18] = 4'b1100;\
game_grid[26][19] = 4'b1100;\
game_grid[26][20] = 4'b1100;\
game_grid[26][21] = 4'b1100;\
game_grid[26][22] = 4'b1100;\
game_grid[26][23] = 4'b1100;\
game_grid[26][24] = 4'b1100;\
game_grid[26][25] = 4'b1100;\
game_grid[26][26] = 4'b1100;\
game_grid[26][27] = 4'b1100;\
game_grid[26][28] = 4'b1100;\
game_grid[26][29] = 4'b1100;\
game_grid[27][0] = 4'b1100;\
game_grid[27][1] = 4'b1100;\
game_grid[27][2] = 4'b1100;\
game_grid[27][3] = 4'b1100;\
game_grid[27][4] = 4'b1100;\
game_grid[27][5] = 4'b1100;\
game_grid[27][6] = 4'b1100;\
game_grid[27][7] = 4'b1100;\
game_grid[27][8] = 4'b1100;\
game_grid[27][9] = 4'b1100;\
game_grid[27][10] = 4'b1100;\
game_grid[27][11] = 4'b1100;\
game_grid[27][12] = 4'b1100;\
game_grid[27][13] = 4'b1100;\
game_grid[27][14] = 4'b1100;\
game_grid[27][15] = 4'b1100;\
game_grid[27][16] = 4'b1100;\
game_grid[27][17] = 4'b1100;\
game_grid[27][18] = 4'b1100;\
game_grid[27][19] = 4'b1100;\
game_grid[27][20] = 4'b1100;\
game_grid[27][21] = 4'b1100;\
game_grid[27][22] = 4'b1100;\
game_grid[27][23] = 4'b1100;\
game_grid[27][24] = 4'b1100;\
game_grid[27][25] = 4'b1100;\
game_grid[27][26] = 4'b1100;\
game_grid[27][27] = 4'b1100;\
game_grid[27][28] = 4'b1100;\
game_grid[27][29] = 4'b1100;\
game_grid[28][0] = 4'b1100;\
game_grid[28][1] = 4'b1100;\
game_grid[28][2] = 4'b1100;\
game_grid[28][3] = 4'b1100;\
game_grid[28][4] = 4'b1100;\
game_grid[28][5] = 4'b1100;\
game_grid[28][6] = 4'b1100;\
game_grid[28][7] = 4'b1100;\
game_grid[28][8] = 4'b1100;\
game_grid[28][9] = 4'b1100;\
game_grid[28][10] = 4'b1100;\
game_grid[28][11] = 4'b1100;\
game_grid[28][12] = 4'b1100;\
game_grid[28][13] = 4'b1100;\
game_grid[28][14] = 4'b1100;\
game_grid[28][15] = 4'b1100;\
game_grid[28][16] = 4'b1100;\
game_grid[28][17] = 4'b1100;\
game_grid[28][18] = 4'b1100;\
game_grid[28][19] = 4'b1100;\
game_grid[28][20] = 4'b1100;\
game_grid[28][21] = 4'b1100;\
game_grid[28][22] = 4'b1100;\
game_grid[28][23] = 4'b1100;\
game_grid[28][24] = 4'b1100;\
game_grid[28][25] = 4'b1100;\
game_grid[28][26] = 4'b1100;\
game_grid[28][27] = 4'b1100;\
game_grid[28][28] = 4'b1100;\
game_grid[28][29] = 4'b1100;\
game_grid[29][0] = 4'b1100;\
game_grid[29][1] = 4'b1100;\
game_grid[29][2] = 4'b1100;\
game_grid[29][3] = 4'b1100;\
game_grid[29][4] = 4'b1100;\
game_grid[29][5] = 4'b1100;\
game_grid[29][6] = 4'b1100;\
game_grid[29][7] = 4'b1100;\
game_grid[29][8] = 4'b1100;\
game_grid[29][9] = 4'b1100;\
game_grid[29][10] = 4'b1100;\
game_grid[29][11] = 4'b1100;\
game_grid[29][12] = 4'b1100;\
game_grid[29][13] = 4'b1100;\
game_grid[29][14] = 4'b1100;\
game_grid[29][15] = 4'b1100;\
game_grid[29][16] = 4'b1100;\
game_grid[29][17] = 4'b1100;\
game_grid[29][18] = 4'b1100;\
game_grid[29][19] = 4'b1100;\
game_grid[29][20] = 4'b1100;\
game_grid[29][21] = 4'b1100;\
game_grid[29][22] = 4'b1100;\
game_grid[29][23] = 4'b1100;\
game_grid[29][24] = 4'b1100;\
game_grid[29][25] = 4'b1100;\
game_grid[29][26] = 4'b1100;\
game_grid[29][27] = 4'b1100;\
game_grid[29][28] = 4'b1100;\
game_grid[29][29] = 4'b1100;\
game_grid[30][0] = 4'b1100;\
game_grid[30][1] = 4'b1100;\
game_grid[30][2] = 4'b1100;\
game_grid[30][3] = 4'b1100;\
game_grid[30][4] = 4'b1100;\
game_grid[30][5] = 4'b1100;\
game_grid[30][6] = 4'b1100;\
game_grid[30][7] = 4'b1100;\
game_grid[30][8] = 4'b1100;\
game_grid[30][9] = 4'b1100;\
game_grid[30][10] = 4'b1100;\
game_grid[30][11] = 4'b1100;\
game_grid[30][12] = 4'b1100;\
game_grid[30][13] = 4'b1100;\
game_grid[30][14] = 4'b1100;\
game_grid[30][15] = 4'b1100;\
game_grid[30][16] = 4'b1100;\
game_grid[30][17] = 4'b1100;\
game_grid[30][18] = 4'b1100;\
game_grid[30][19] = 4'b1100;\
game_grid[30][20] = 4'b1100;\
game_grid[30][21] = 4'b1100;\
game_grid[30][22] = 4'b1100;\
game_grid[30][23] = 4'b1100;\
game_grid[30][24] = 4'b1100;\
game_grid[30][25] = 4'b1100;\
game_grid[30][26] = 4'b1100;\
game_grid[30][27] = 4'b1100;\
game_grid[30][28] = 4'b1100;\
game_grid[30][29] = 4'b1100;\
game_grid[31][0] = 4'b1100;\
game_grid[31][1] = 4'b1100;\
game_grid[31][2] = 4'b1100;\
game_grid[31][3] = 4'b1100;\
game_grid[31][4] = 4'b1100;\
game_grid[31][5] = 4'b1100;\
game_grid[31][6] = 4'b1100;\
game_grid[31][7] = 4'b1100;\
game_grid[31][8] = 4'b1100;\
game_grid[31][9] = 4'b1100;\
game_grid[31][10] = 4'b1100;\
game_grid[31][11] = 4'b1100;\
game_grid[31][12] = 4'b1100;\
game_grid[31][13] = 4'b1100;\
game_grid[31][14] = 4'b1100;\
game_grid[31][15] = 4'b1100;\
game_grid[31][16] = 4'b1100;\
game_grid[31][17] = 4'b1100;\
game_grid[31][18] = 4'b1100;\
game_grid[31][19] = 4'b1100;\
game_grid[31][20] = 4'b1100;\
game_grid[31][21] = 4'b1100;\
game_grid[31][22] = 4'b1100;\
game_grid[31][23] = 4'b1100;\
game_grid[31][24] = 4'b1100;\
game_grid[31][25] = 4'b1100;\
game_grid[31][26] = 4'b1100;\
game_grid[31][27] = 4'b1100;\
game_grid[31][28] = 4'b1100;\
game_grid[31][29] = 4'b1100;\
game_grid[32][0] = 4'b1100;\
game_grid[32][1] = 4'b1100;\
game_grid[32][2] = 4'b1100;\
game_grid[32][3] = 4'b1100;\
game_grid[32][4] = 4'b1100;\
game_grid[32][5] = 4'b1100;\
game_grid[32][6] = 4'b1100;\
game_grid[32][7] = 4'b1100;\
game_grid[32][8] = 4'b1100;\
game_grid[32][9] = 4'b1100;\
game_grid[32][10] = 4'b1100;\
game_grid[32][11] = 4'b1100;\
game_grid[32][12] = 4'b1100;\
game_grid[32][13] = 4'b1100;\
game_grid[32][14] = 4'b1100;\
game_grid[32][15] = 4'b1100;\
game_grid[32][16] = 4'b1100;\
game_grid[32][17] = 4'b1100;\
game_grid[32][18] = 4'b1100;\
game_grid[32][19] = 4'b1100;\
game_grid[32][20] = 4'b1100;\
game_grid[32][21] = 4'b1100;\
game_grid[32][22] = 4'b1100;\
game_grid[32][23] = 4'b1100;\
game_grid[32][24] = 4'b1100;\
game_grid[32][25] = 4'b1100;\
game_grid[32][26] = 4'b1100;\
game_grid[32][27] = 4'b1100;\
game_grid[32][28] = 4'b1100;\
game_grid[32][29] = 4'b1100;\
game_grid[33][0] = 4'b1100;\
game_grid[33][1] = 4'b1100;\
game_grid[33][2] = 4'b1100;\
game_grid[33][3] = 4'b1100;\
game_grid[33][4] = 4'b1100;\
game_grid[33][5] = 4'b1100;\
game_grid[33][6] = 4'b1100;\
game_grid[33][7] = 4'b1100;\
game_grid[33][8] = 4'b1100;\
game_grid[33][9] = 4'b1100;\
game_grid[33][10] = 4'b1100;\
game_grid[33][11] = 4'b1100;\
game_grid[33][12] = 4'b1100;\
game_grid[33][13] = 4'b1100;\
game_grid[33][14] = 4'b1100;\
game_grid[33][15] = 4'b1100;\
game_grid[33][16] = 4'b1100;\
game_grid[33][17] = 4'b1100;\
game_grid[33][18] = 4'b1100;\
game_grid[33][19] = 4'b1100;\
game_grid[33][20] = 4'b1100;\
game_grid[33][21] = 4'b1100;\
game_grid[33][22] = 4'b1100;\
game_grid[33][23] = 4'b1100;\
game_grid[33][24] = 4'b1100;\
game_grid[33][25] = 4'b1100;\
game_grid[33][26] = 4'b1100;\
game_grid[33][27] = 4'b1100;\
game_grid[33][28] = 4'b1100;\
game_grid[33][29] = 4'b1100;\
game_grid[34][0] = 4'b1100;\
game_grid[34][1] = 4'b1100;\
game_grid[34][2] = 4'b1100;\
game_grid[34][3] = 4'b1100;\
game_grid[34][4] = 4'b1100;\
game_grid[34][5] = 4'b1100;\
game_grid[34][6] = 4'b1100;\
game_grid[34][7] = 4'b1100;\
game_grid[34][8] = 4'b1100;\
game_grid[34][9] = {`ENT_APPLE, 2'b00};\
game_grid[34][10] = 4'b1100;\
game_grid[34][11] = 4'b1100;\
game_grid[34][12] = 4'b1100;\
game_grid[34][13] = 4'b1100;\
game_grid[34][14] = 4'b1100;\
game_grid[34][15] = 4'b1100;\
game_grid[34][16] = 4'b1100;\
game_grid[34][17] = 4'b1100;\
game_grid[34][18] = 4'b1100;\
game_grid[34][19] = 4'b1100;\
game_grid[34][20] = 4'b1100;\
game_grid[34][21] = 4'b1100;\
game_grid[34][22] = 4'b1100;\
game_grid[34][23] = 4'b1100;\
game_grid[34][24] = 4'b1100;\
game_grid[34][25] = 4'b1100;\
game_grid[34][26] = 4'b1100;\
game_grid[34][27] = 4'b1100;\
game_grid[34][28] = 4'b1100;\
game_grid[34][29] = 4'b1100;\
game_grid[35][0] = 4'b1100;\
game_grid[35][1] = 4'b1100;\
game_grid[35][2] = 4'b1100;\
game_grid[35][3] = 4'b1100;\
game_grid[35][4] = 4'b1100;\
game_grid[35][5] = 4'b1100;\
game_grid[35][6] = 4'b1100;\
game_grid[35][7] = 4'b1100;\
game_grid[35][8] = 4'b1100;\
game_grid[35][9] = 4'b1100;\
game_grid[35][10] = 4'b1100;\
game_grid[35][11] = 4'b1100;\
game_grid[35][12] = 4'b1100;\
game_grid[35][13] = 4'b1100;\
game_grid[35][14] = 4'b1100;\
game_grid[35][15] = 4'b1100;\
game_grid[35][16] = 4'b1100;\
game_grid[35][17] = 4'b1100;\
game_grid[35][18] = 4'b1100;\
game_grid[35][19] = 4'b1100;\
game_grid[35][20] = 4'b1100;\
game_grid[35][21] = 4'b1100;\
game_grid[35][22] = 4'b1100;\
game_grid[35][23] = 4'b1100;\
game_grid[35][24] = 4'b1100;\
game_grid[35][25] = 4'b1100;\
game_grid[35][26] = 4'b1100;\
game_grid[35][27] = 4'b1100;\
game_grid[35][28] = 4'b1100;\
game_grid[35][29] = 4'b1100;\
game_grid[36][0] = 4'b1100;\
game_grid[36][1] = 4'b1100;\
game_grid[36][2] = 4'b1100;\
game_grid[36][3] = 4'b1100;\
game_grid[36][4] = 4'b1100;\
game_grid[36][5] = 4'b1100;\
game_grid[36][6] = 4'b1100;\
game_grid[36][7] = 4'b1100;\
game_grid[36][8] = 4'b1100;\
game_grid[36][9] = 4'b1100;\
game_grid[36][10] = 4'b1100;\
game_grid[36][11] = 4'b1100;\
game_grid[36][12] = 4'b1100;\
game_grid[36][13] = 4'b1100;\
game_grid[36][14] = 4'b1100;\
game_grid[36][15] = 4'b1100;\
game_grid[36][16] = 4'b1100;\
game_grid[36][17] = 4'b1100;\
game_grid[36][18] = 4'b1100;\
game_grid[36][19] = 4'b1100;\
game_grid[36][20] = 4'b1100;\
game_grid[36][21] = 4'b1100;\
game_grid[36][22] = 4'b1100;\
game_grid[36][23] = 4'b1100;\
game_grid[36][24] = 4'b1100;\
game_grid[36][25] = 4'b1100;\
game_grid[36][26] = 4'b1100;\
game_grid[36][27] = 4'b1100;\
game_grid[36][28] = 4'b1100;\
game_grid[36][29] = 4'b1100;\
game_grid[37][0] = 4'b1100;\
game_grid[37][1] = 4'b1100;\
game_grid[37][2] = 4'b1100;\
game_grid[37][3] = 4'b1100;\
game_grid[37][4] = 4'b1100;\
game_grid[37][5] = 4'b1100;\
game_grid[37][6] = 4'b1100;\
game_grid[37][7] = 4'b1100;\
game_grid[37][8] = 4'b1100;\
game_grid[37][9] = 4'b1100;\
game_grid[37][10] = 4'b1100;\
game_grid[37][11] = 4'b1100;\
game_grid[37][12] = 4'b1100;\
game_grid[37][13] = 4'b1100;\
game_grid[37][14] = 4'b1100;\
game_grid[37][15] = 4'b1100;\
game_grid[37][16] = 4'b1100;\
game_grid[37][17] = 4'b1100;\
game_grid[37][18] = 4'b1100;\
game_grid[37][19] = 4'b1100;\
game_grid[37][20] = 4'b1100;\
game_grid[37][21] = 4'b1100;\
game_grid[37][22] = 4'b1100;\
game_grid[37][23] = 4'b1100;\
game_grid[37][24] = 4'b1100;\
game_grid[37][25] = 4'b1100;\
game_grid[37][26] = 4'b1100;\
game_grid[37][27] = 4'b1100;\
game_grid[37][28] = 4'b1100;\
game_grid[37][29] = 4'b1100;\
game_grid[38][0] = 4'b1100;\
game_grid[38][1] = 4'b1100;\
game_grid[38][2] = 4'b1100;\
game_grid[38][3] = 4'b1100;\
game_grid[38][4] = 4'b1100;\
game_grid[38][5] = 4'b1100;\
game_grid[38][6] = 4'b1100;\
game_grid[38][7] = 4'b1100;\
game_grid[38][8] = 4'b1100;\
game_grid[38][9] = 4'b1100;\
game_grid[38][10] = 4'b1100;\
game_grid[38][11] = 4'b1100;\
game_grid[38][12] = 4'b1100;\
game_grid[38][13] = 4'b1100;\
game_grid[38][14] = 4'b1100;\
game_grid[38][15] = 4'b1100;\
game_grid[38][16] = 4'b1100;\
game_grid[38][17] = 4'b1100;\
game_grid[38][18] = 4'b1100;\
game_grid[38][19] = 4'b1100;\
game_grid[38][20] = 4'b1100;\
game_grid[38][21] = 4'b1100;\
game_grid[38][22] = 4'b1100;\
game_grid[38][23] = 4'b1100;\
game_grid[38][24] = 4'b1100;\
game_grid[38][25] = 4'b1100;\
game_grid[38][26] = 4'b1100;\
game_grid[38][27] = 4'b1100;\
game_grid[38][28] = 4'b1100;\
game_grid[38][29] = 4'b1100;\
game_grid[39][0] = 4'b1100;\
game_grid[39][1] = 4'b1100;\
game_grid[39][2] = 4'b1100;\
game_grid[39][3] = 4'b1100;\
game_grid[39][4] = 4'b1100;\
game_grid[39][5] = 4'b1100;\
game_grid[39][6] = 4'b1100;\
game_grid[39][7] = 4'b1100;\
game_grid[39][8] = 4'b1100;\
game_grid[39][9] = 4'b1100;\
game_grid[39][10] = 4'b1100;\
game_grid[39][11] = 4'b1100;\
game_grid[39][12] = 4'b1100;\
game_grid[39][13] = 4'b1100;\
game_grid[39][14] = 4'b1100;\
game_grid[39][15] = 4'b1100;\
game_grid[39][16] = 4'b1100;\
game_grid[39][17] = 4'b1100;\
game_grid[39][18] = 4'b1100;\
game_grid[39][19] = 4'b1100;\
game_grid[39][20] = 4'b1100;\
game_grid[39][21] = 4'b1100;\
game_grid[39][22] = 4'b1100;\
game_grid[39][23] = 4'b1100;\
game_grid[39][24] = 4'b1100;\
game_grid[39][25] = 4'b1100;\
game_grid[39][26] = 4'b1100;\
game_grid[39][27] = 4'b1100;\
game_grid[39][28] = 4'b1100;\
game_grid[39][29] = 4'b1100;\

`endif // init_vh
